


module  c6 ( input Reset, frame_clk, input [7:0] keycode,
               output [9:0]  C6X, C6Y);
    
       
    assign C6X = 450;
   
    assign C6Y = 300;
    

endmodule
