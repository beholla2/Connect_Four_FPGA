


module  b2 ( input Reset, frame_clk, input [7:0] keycode,
               output [9:0]  B2X, B2Y);
    
       
    assign B2X = 150;
   
    assign B2Y = 375;
    

endmodule
