


module  e6 ( input Reset, frame_clk, input [7:0] keycode,
               output [9:0]  E6X, E6Y);
    
       
    assign E6X = 450;
   
    assign E6Y = 150;
    

endmodule
