


module  e2 ( input Reset, frame_clk, input [7:0] keycode,
               output [9:0]  E2X, E2Y);
    
       
    assign E2X = 150;
   
    assign E2Y = 150;
    

endmodule
