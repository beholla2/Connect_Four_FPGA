


module  e4 ( input Reset, frame_clk, input [7:0] keycode,
               output [9:0]  E4X, E4Y);
    
       
    assign E4X = 300;
   
    assign E4Y = 150;
    

endmodule
