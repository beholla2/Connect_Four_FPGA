


module  d6 ( input Reset, frame_clk, input [7:0] keycode,
               output [9:0]  D6X, D6Y);
    
       
    assign D6X = 450;
   
    assign D6Y = 225;
    

endmodule
