// Module for drawing the board

module  f5 ( input Reset, frame_clk, input [7:0] keycode,
               output [9:0]  F5X, F5Y);
    
       
    assign F5X = 375;
   
    assign F5Y = 75;
    

endmodule
