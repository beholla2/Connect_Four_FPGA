


module  e1 ( input Reset, frame_clk, input [7:0] keycode,
               output [9:0]  E1X, E1Y);
    
       
    assign E1X = 75;
   
    assign E1Y = 150;
    

endmodule
