


module  c1 ( input Reset, frame_clk, input [7:0] keycode,
               output [9:0]  C1X, C1Y);
    
       
    assign C1X = 75;
   
    assign C1Y = 300;
    

endmodule
