


module  b6 ( input Reset, frame_clk, input [7:0] keycode,
               output [9:0]  B6X, B6Y);
    
       
    assign B6X = 450;
   
    assign B6Y = 375;
    

endmodule
