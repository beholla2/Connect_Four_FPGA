


module  c2 ( input Reset, frame_clk, input [7:0] keycode,
               output [9:0]  C2X, C2Y);
    
       
    assign C2X = 150;
   
    assign C2Y = 300;
    

endmodule
