


module  c3 ( input Reset, frame_clk, input [7:0] keycode,
               output [9:0]  C3X, C3Y);
    
       
    assign C3X = 225;
   
    assign C3Y = 300;
    

endmodule
