


module  b3 ( input Reset, frame_clk, input [7:0] keycode,
               output [9:0]  B3X, B3Y);
    
       
    assign B3X = 225;
   
    assign B3Y = 375;
    

endmodule
