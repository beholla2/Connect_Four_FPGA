


module  c7 ( input Reset, frame_clk, input [7:0] keycode,
               output [9:0]  C7X, C7Y);
    
       
    assign C7X = 525;
   
    assign C7Y = 300;
    

endmodule
