


module  c5 ( input Reset, frame_clk, input [7:0] keycode,
               output [9:0]  C5X, C5Y);
    
       
    assign C5X = 375;
   
    assign C5Y = 300;
    

endmodule
