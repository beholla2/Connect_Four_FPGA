


module  e7 ( input Reset, frame_clk, input [7:0] keycode,
               output [9:0]  E7X, E7Y);
    
       
    assign E7X = 525;
   
    assign E7Y = 150;
    

endmodule
