


module  b4 ( input Reset, frame_clk, input [7:0] keycode,
               output [9:0]  B4X, B4Y);
    
       
    assign B4X = 300;
   
    assign B4Y = 375;
    

endmodule
