


module  d2 ( input Reset, frame_clk, input [7:0] keycode,
               output [9:0]  D2X, D2Y);
    
       
    assign D2X = 150;
   
    assign D2Y = 225;
    

endmodule
