


module  d1 ( input Reset, frame_clk, input [7:0] keycode,
               output [9:0]  D1X, D1Y);
    
       
    assign D1X = 75;
   
    assign D1Y = 225;
    

endmodule
