


module  d7 ( input Reset, frame_clk, input [7:0] keycode,
               output [9:0]  D7X, D7Y);
    
       
    assign D7X = 525;
   
    assign D7Y = 225;
    

endmodule
