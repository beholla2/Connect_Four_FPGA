


module  c4 ( input Reset, frame_clk, input [7:0] keycode,
               output [9:0]  C4X, C4Y);
    
       
    assign C4X = 300;
   
    assign C4Y = 300;
    

endmodule
