


module  b5 ( input Reset, frame_clk, input [7:0] keycode,
               output [9:0]  B5X, B5Y);
    
       
    assign B5X = 375;
   
    assign B5Y = 375;
    

endmodule
