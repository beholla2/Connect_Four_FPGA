


module  e5 ( input Reset, frame_clk, input [7:0] keycode,
               output [9:0]  E5X, E5Y);
    
       
    assign E5X = 375;
   
    assign E5Y = 150;
    

endmodule
