


module  e3 ( input Reset, frame_clk, input [7:0] keycode,
               output [9:0]  E3X, E3Y);
    
       
    assign E3X = 225;
   
    assign E3Y = 150;
    

endmodule
