// Module for drawing the board

module  f6 ( input Reset, frame_clk, input [7:0] keycode,
               output [9:0]  F6X, F6Y);
    
       
    assign F6X = 450;
   
    assign F6Y = 75;
    

endmodule
