


module  d3 ( input Reset, frame_clk, input [7:0] keycode,
               output [9:0]  D3X, D3Y);
    
       
    assign D3X = 225;
   
    assign D3Y = 225;
    

endmodule
