// Module for drawing the board

module  f7 ( input Reset, frame_clk, input [7:0] keycode,
               output [9:0]  F7X, F7Y);
    
       
    assign F7X = 525;
   
    assign F7Y = 75;
    

endmodule
