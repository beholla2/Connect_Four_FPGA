


module  b1 ( input Reset, frame_clk, input [7:0] keycode,
               output [9:0]  B1X, B1Y);
    
       
    assign B1X = 75;
   
    assign B1Y = 375;
    

endmodule
