


module  b7 ( input Reset, frame_clk, input [7:0] keycode,
               output [9:0]  B7X, B7Y);
    
       
    assign B7X = 525;
   
    assign B7Y = 375;
    

endmodule
