


module  d4 ( input Reset, frame_clk, input [7:0] keycode,
               output [9:0]  D4X, D4Y);
    
       
    assign D4X = 300;
   
    assign D4Y = 225;
    

endmodule
