


module  d5 ( input Reset, frame_clk, input [7:0] keycode,
               output [9:0]  D5X, D5Y);
    
       
    assign D5X = 375;
   
    assign D5Y = 225;
    

endmodule
